library verilog;
use verilog.vl_types.all;
entity Completo_vlg_vec_tst is
end Completo_vlg_vec_tst;
