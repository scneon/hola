-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Sun Dec 11 20:34:38 2022

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ProyectoTyDD2 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        N : IN STD_LOGIC := '0';
        Z2 : OUT STD_LOGIC;
        Z1 : OUT STD_LOGIC;
        Z0 : OUT STD_LOGIC
    );
END ProyectoTyDD2;

ARCHITECTURE BEHAVIOR OF ProyectoTyDD2 IS
    TYPE type_fstate IS (A_000,B_100,C_110,D_010,E_111,F_101,G_011,H_001,I_110,J_111,K_100,L_101,M_010,N_011,O_001,P_000);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,N)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= A_000;
            Z2 <= '0';
            Z1 <= '0';
            Z0 <= '0';
        ELSE
            Z2 <= '0';
            Z1 <= '0';
            Z0 <= '0';
            CASE fstate IS
                WHEN A_000 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= A_000;
                    ELSIF ((N = '0')) THEN
                        reg_fstate <= B_100;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= A_000;
                    END IF;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z2 <= '0';
                WHEN B_100 =>
                    IF ((N = '0')) THEN
                        reg_fstate <= C_110;
                    ELSIF ((N = '1')) THEN
                        reg_fstate <= D_010;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= B_100;
                    END IF;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z2 <= '1';
                WHEN C_110 =>
                    IF ((N = '0')) THEN
                        reg_fstate <= E_111;
                    ELSIF ((N = '1')) THEN
                        reg_fstate <= F_101;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= C_110;
                    END IF;

                    Z0 <= '0';

                    Z1 <= '1';

                    Z2 <= '1';
                WHEN D_010 =>
                    IF ((N = '0')) THEN
                        reg_fstate <= G_011;
                    ELSIF ((N = '1')) THEN
                        reg_fstate <= H_001;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= D_010;
                    END IF;

                    Z0 <= '0';

                    Z1 <= '1';

                    Z2 <= '0';
                WHEN E_111 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= I_110;
                    ELSIF ((N = '0')) THEN
                        reg_fstate <= J_111;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= E_111;
                    END IF;

                    Z0 <= '1';

                    Z1 <= '1';

                    Z2 <= '1';
                WHEN F_101 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= K_100;
                    ELSIF ((N = '0')) THEN
                        reg_fstate <= L_101;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= F_101;
                    END IF;

                    Z0 <= '1';

                    Z1 <= '0';

                    Z2 <= '1';
                WHEN G_011 =>
                    IF ((N = '1')) THEN
                        reg_fstate <= M_010;
                    ELSIF ((N = '0')) THEN
                        reg_fstate <= N_011;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= G_011;
                    END IF;

                    Z0 <= '1';

                    Z1 <= '1';

                    Z2 <= '0';
                WHEN H_001 =>
                    IF ((N = '0')) THEN
                        reg_fstate <= O_001;
                    ELSIF ((N = '1')) THEN
                        reg_fstate <= P_000;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= H_001;
                    END IF;

                    Z0 <= '1';

                    Z1 <= '0';

                    Z2 <= '0';
                WHEN I_110 =>
                    reg_fstate <= I_110;

                    Z0 <= '0';

                    Z1 <= '1';

                    Z2 <= '1';
                WHEN J_111 =>
                    reg_fstate <= J_111;

                    Z0 <= '1';

                    Z1 <= '1';

                    Z2 <= '1';
                WHEN K_100 =>
                    reg_fstate <= K_100;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z2 <= '1';
                WHEN L_101 =>
                    reg_fstate <= L_101;

                    Z0 <= '1';

                    Z1 <= '0';

                    Z2 <= '1';
                WHEN M_010 =>
                    reg_fstate <= M_010;

                    Z0 <= '0';

                    Z1 <= '1';

                    Z2 <= '0';
                WHEN N_011 =>
                    reg_fstate <= N_011;

                    Z0 <= '1';

                    Z1 <= '1';

                    Z2 <= '0';
                WHEN O_001 =>
                    reg_fstate <= O_001;

                    Z0 <= '1';

                    Z1 <= '0';

                    Z2 <= '0';
                WHEN P_000 =>
                    reg_fstate <= P_000;

                    Z0 <= '0';

                    Z1 <= '0';

                    Z2 <= '0';
                WHEN OTHERS => 
                    Z2 <= 'X';
                    Z1 <= 'X';
                    Z0 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
